`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/18/2020 08:42:58 PM
// Design Name: 
// Module Name: all2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


// -------------------------------------------------------------
// 
// File Name: hdlsrc/test2/test2.v
// Created: 2020-03-18 16:04:18
// 
// Generated by MATLAB 9.7 and HDL Coder 3.15
// 
// 
// -- -------------------------------------------------------------
// -- Rate and Clocking Details
// -- -------------------------------------------------------------
// Model base rate: 1e-08
// Target subsystem base rate: 1e-08
// 
// -------------------------------------------------------------


// -------------------------------------------------------------
// 
// Module: test2
// Source Path: test2
// Hierarchy Level: 0
// 
// -------------------------------------------------------------

`timescale 1 ns / 1 ns

module all2
          (clk,
           resetn,
           //clk_enable,
           SW,
           PDM,
           JA,
           AUD_SD);


  input   clk;
  input   resetn;
  //input   clk_enable;
  input   [15:0] SW;
  output  PDM;
  output  [4:1] JA;
  output  AUD_SD;
  assign AUD_SD = 1;
  wire   PDM_mid;

  wire signed [19:0] HDL_DUT_out2;  // sfix20_En18
  wire signed [19:0] HDL_DUT_out3;  // sfix20_En18
  wire signed [19:0] HDL_DUT_out4;  // sfix20_En18
  wire signed [19:0] HDL_DUT_out5;  // sfix20_En18
  wire signed [23:0] HDL_DUT_out6;  // sfix24_En14
  wire signed [23:0] HDL_DUT_out7;  // sfix24_En14

  // Note: This model is configured with 'hdlsetup'
  // 
  // Add your design targeted for ASIC/FPGA inside HDL_DUT and then run the following command:
  // makehdl('HDL_DUT')
  // 
  // Copyright 2015-2016 The MathWorks, Inc.

  assign JA[1] = PDM;
  assign JA[2] = PDM;
  assign JA[3] = PDM;
  assign JA[4] = PDM;
  //assign JA[5] = PDM;
  //assign JA[6] = PDM;
//  assign JA[7] = PDM;
//  assign JA[8] = PDM;
//  assign JA[9] = PDM;
//  assign JA[10]= PDM;
  
  HDL_DUT u_HDL_DUT (.clk(clk),
                     .reset(~resetn),
                     .clk_enable(1),
                     .ce_out(),
                     .Input1(SW[0]),
                     .Input2(SW[1]),
                     .Input3(SW[2]),
                     .Input4(SW[3]),
                     .run_drum(SW[4]),
                     //.rst_drum(SW[5]),
                     .out1(PDM_mid),
                     .out(HDL_DUT_out2),  // sfix20_En18
                     .out2(HDL_DUT_out3),  // sfix20_En18
                     .out3(HDL_DUT_out4),  // sfix20_En18
                     .out4(HDL_DUT_out5),  // sfix20_En18
                     .Integrator(HDL_DUT_out6),  // sfix24_En14
                     .Unmodulated(HDL_DUT_out7)  // sfix24_En14
                     );
    assign PDM = PDM_mid & (SW[0] | SW[1] | SW[2] | SW[3] | SW[4]);
endmodule  // test2

